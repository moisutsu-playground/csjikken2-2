/******************/
/* signext16_32.v */
/******************/

//            +----+
//  sign_ext->|    |
// a16[15:0]->|    |->y32[31:0]
//            +----+

module signext16_32 (sign_ext, a16, y32);  // 入出力ポート
  input      sign_ext;          // 入力 1-bit
  input   [15:0]  a16;          // 入力 16-bit
  output  [31:0]  y32;          // 出力 32-bit

  //Body
  //符号拡張
  assign y32 = (sign_ext == 1'b1) ?
               {a16[15], a16[15], a16[15], a16[15],
                a16[15], a16[15], a16[15], a16[15],
                a16[15], a16[15], a16[15], a16[15],
                a16[15], a16[15], a16[15], a16[15],
                a16[15:0]}
               : {16'h0000, a16[15:0]};
endmodule
