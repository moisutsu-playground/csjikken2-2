library verilog;
use verilog.vl_types.all;
entity test_cpu is
end test_cpu;
